library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.HermesPackage.all;

package TablePackage is

constant NREG : integer := 4;
constant MEMORY_SIZE : integer := NREG;
constant NBITS : integer := 2;
constant CELL_SIZE : integer := 2*NPORT+4*NBITS;

subtype cell is std_logic_vector(CELL_SIZE-1 downto 0);
type memory is array (0 to MEMORY_SIZE-1) of cell;
type tables is array (0 to NROT-1) of memory;

constant TAB: tables :=(
 -- Router 0.0
(("100000001001100100"),
("100000100111100001"),
("000000000000000000"),
("000000000000000000")
),
 -- Router 0.1
(("000000100110100001"),
("000000010111100100"),
("000000000000001000"),
("000000000000000000")
),
 -- Router 0.2
(("000000011001100100"),
("000000000000101000"),
("000000100111100001"),
("000000000000000000")
),
 -- Router 0.3
(("100000000001001000"),
("100000100111100001"),
("000000000000000000"),
("000000000000000000")
),
 -- Router 1.0
(("000000000000000010"),
("000000001011100100"),
("000001000111100001"),
("000000000000000000")
),
 -- Router 1.1
(("000000000010001000"),
("000000000000100010"),
("000001000110100001"),
("000000010111100100")
),
 -- Router 1.2
(("000000100010101000"),
("000000011011100100"),
("000000000001000010"),
("000001000111100001")
),
 -- Router 1.3
(("000000011001100010"),
("000000000011001000"),
("000001000111100001"),
("000000000000000000")
),
 -- Router 2.0
(("000000000010000010"),
("000001100111100001"),
("000000001101100100"),
("000000000000000000")
),
 -- Router 2.1
(("000001100110100001"),
("000000000100001000"),
("000000000010100010"),
("000000010111100100")
),
 -- Router 2.2
(("000001000100101000"),
("000001100111000001"),
("000000011111100100"),
("000000000011000010")
),
 -- Router 2.3
(("000000011011100010"),
("000001100111100001"),
("000000000101001000"),
("000000000000000000")
),
 -- Router 3.0
(("000000001111100100"),
("000000000100000010"),
("000000000000000000"),
("000000000000000000")
),
 -- Router 3.1
(("000000000110001000"),
("000000000100100010"),
("000000010111100100"),
("000000000000000000")
),
 -- Router 3.2
(("000001100110101000"),
("000000000100001000"),
("000000011111100100"),
("000000000101000010")
),
 -- Router 3.3
(("000001100111001000"),
("000000000101100010"),
("000000000000000000"),
("000000000000000000")
)
);
end TablePackage;

package body TablePackage is
end TablePackage;
